library verilog;
use verilog.vl_types.all;
entity Main_Decoder_tb is
end Main_Decoder_tb;
