library verilog;
use verilog.vl_types.all;
entity Core_Datapath_tb is
end Core_Datapath_tb;
