library verilog;
use verilog.vl_types.all;
entity Extend_tb is
end Extend_tb;
