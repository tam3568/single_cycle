library verilog;
use verilog.vl_types.all;
entity Instruction_Memory_tb is
end Instruction_Memory_tb;
