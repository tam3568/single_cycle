library verilog;
use verilog.vl_types.all;
entity PC_Plus_4_tb is
end PC_Plus_4_tb;
