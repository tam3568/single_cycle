library verilog;
use verilog.vl_types.all;
entity Result_Mux_tb is
end Result_Mux_tb;
