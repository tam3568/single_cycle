library verilog;
use verilog.vl_types.all;
entity Single_Cycle_TB is
end Single_Cycle_TB;
