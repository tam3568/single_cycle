library verilog;
use verilog.vl_types.all;
entity Register_File_tb is
end Register_File_tb;
