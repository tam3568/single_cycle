library verilog;
use verilog.vl_types.all;
entity ALU_Decoder_tb is
end ALU_Decoder_tb;
