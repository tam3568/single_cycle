library verilog;
use verilog.vl_types.all;
entity PC_Target_tb is
end PC_Target_tb;
