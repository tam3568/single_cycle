library verilog;
use verilog.vl_types.all;
entity ALU_Mux_tb is
end ALU_Mux_tb;
