library verilog;
use verilog.vl_types.all;
entity PC_Mux_tb is
end PC_Mux_tb;
